module digital_design_lab1_problem3
	#(parameter n = 6)
	(input logic reset, dcrease_btn, output logic isNegative, output logic [n-1:0] value, output logic [6:0] segUnits, segDec, segSign);
	
	
	
	